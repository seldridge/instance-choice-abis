module Baz(output a);
  assign a = 1'h1;
endmodule
