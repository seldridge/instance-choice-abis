module Baz();
  wire a = 1'h1;
endmodule
