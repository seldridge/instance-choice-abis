module Test();

  Foo foo();
  wire a = foo.`ref_Foo_x;

endmodule
