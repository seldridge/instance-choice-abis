module Bar(output a);
  assign a = 1'h0;
endmodule
