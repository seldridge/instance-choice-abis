module Bar();
  wire b = 1'h0;
endmodule
