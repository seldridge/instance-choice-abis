// Defines for probes associated with module `Foo`.

`ifndef __targetref_Foo_x_a
 `define __targetref_Foo_x_a b
`endif

`define ref_Foo_x x.`__targetref_Foo_x_a
